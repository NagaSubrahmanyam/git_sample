4. From working directory to staging area we will use a command called git add <file name>. Then that file removed from untracked files list

1. Without this area we can't able to send only required no of files to local repository.
2. First we will send how many files we want send to local repository those many we can send to Staging area. Form there we can send all the files to local repository.
3. After adding the files to staging area those files will comes under Changes to be committed list.

